module binary_to_hex_7segDecoder ();


endmodule 